/* top-level divider circuit for use in homework 4.
 *
 * Inputs:
 *   Clock  - should be connected to a 50 MHz clock
 *   Resetn - negated reset (resets on 0)
 *   s      - signal to start running
 *   DataA  - numerator/dividend number for division
 *   DataB  - denominator/divisor number for division
 *
 * Outputs:
 *   R     - remainder from division
 *   Q     - quotient from division
 *   Done  - signal circut finished dividing
 *
 * Parameters:
 *   n     - bit-length of input nums
 *   logn  - log base 2 of the bit-length of input nums
 *
 * CHANGE: Removed LA, EB from input ports, should be generated by controller
 */
module divider (Clock, Resetn, s, DataA, DataB, R, Q, Done);
	parameter n = 8, logn = 3;
	input Clock, Resetn, s;
	input [n-1:0] DataA, DataB;
	output [n-1:0] R, Q;
	output logic Done;
	
	logic Cout, z;
	logic [n-1:0] DataR;
	logic [n:0] Sum;
	logic [1:0] y, Y;
	logic [n-1:0] A, B;
	logic [logn-1:0] Count;
	logic EA, Rsel, LR, ER, ER0, LC, EC, R0, LA, EB;
	integer k;

// control circuit

	parameter S1 = 2'b00, S2 = 2'b01, S3 = 2'b10;

	// CHANGE: made pure combinational
	always_comb
	begin: State_table
		case (y)
			S1:	if (s == 0) Y = S1;
				else Y = S2;
			// CHANGE 
			S2:	if (~z) Y = S2;
				else Y = S3;
			S3:	if (s == 1) Y = S3;
				else Y = S1;
			default: Y = 2'bxx;
		endcase
	end

	// CHANGE: made pure sequential
	always_ff @(posedge Clock, negedge Resetn)
	begin: State_flipflops
		if (Resetn == 0)
			y <= S1;
		else
			y <= Y;
	end

	// CHANGE: made pure combinational
	always_comb
	begin: FSM_outputs
		// defaults
		LR = 0; ER = 0; ER0 = 0; LC = 0; EC = 0; EA = 0; LA = 0; EB = 0;	
		Rsel = 0; Done = 0;
		case (y)
			S1:	begin
					LC = 1; ER = 1;
					if (s == 0)
					begin
						LR = 1; ER0 = 0; LA = 1; EB = 1;
					end
					else
					begin
						LR = 0; EA = 1; ER0 = 1;
					end
				end
			S2:	begin
					Rsel = 1; ER = 1; ER0 = 1; EA = 1;
					if (Cout) LR = 1;
					else LR = 0;
					if (~z) EC = 1;
					else EC = 0;
				end
			S3:	Done = 1;
		endcase
	end

//datapath circuit

	regne RegB (DataB, Clock, Resetn, EB, B);
		defparam RegB.n = n;
		
	shiftlne ShiftR (DataR, LR, ER, R0, Clock, R);
		defparam ShiftR.n = n;
		
	muxdff FF_R0 (1'b0, A[n-1], ER0, Clock, R0);
	
	shiftlne ShiftA (DataA, LA, EA, Cout, Clock, A);
		defparam ShiftA.n = n;
		
	assign Q = A;
	
	// CHANGE: Changed load value for counter from 0 -> n-1
	downcount Counter ({logn{1'b1}}, Clock, EC, LC, Count);
		defparam Counter.n = logn;

	assign z = (Count == {logn{1'b0}});

	assign Sum = {1'b0, R[n-2:0], R0} + {1'b0, ~B - '1};
	assign Cout = Sum[n];
	
	// define the n 2-to-1 multiplexers
	assign DataR = Rsel ? Sum : 0;

endmodule

module divider_testbench();
	parameter n = 8;

	logic Clock, Resetn, s, Done, clk;
	logic [n-1:0] DataA, DataB, R, Q;
	
	assign Clock = clk;
	
	divider #(.n(n), .logn(3)) dut (.*);
	
	parameter CLOCK_PERIOD = 100;
	initial begin
		clk <= 0;
		forever #(CLOCK_PERIOD / 2) clk <= ~clk;
	end
	
	initial begin
		integer i;
		
		@(posedge clk) Resetn <= 1'b0; s <= 1'b0; DataA <= 8'd11; DataB <= 4'd2;
		@(posedge clk) Resetn <= 1'b1;
		@(posedge clk);
		@(posedge clk);
		@(posedge clk);
		@(posedge clk); s <= 1'b1;
		
		for (i = 0; i < 10; i++) begin
			@(posedge clk);
		end
		
		@(posedge clk) s <= 1'b0; DataA <= 8'd239; DataB <= 8'd17;
		@(posedge clk);
		@(posedge clk);
		@(posedge clk);
		@(posedge clk); s <= 1'b1;
		for (i = 0; i < 10; i++) begin
			@(posedge clk);
		end
		
		$stop;
	end


endmodule  // divider_testbench

