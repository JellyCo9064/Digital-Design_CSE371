// Code from "FPGA prototyping by SystemVerilog examples" by P. Chu
// Implements a 4-bit sign-and-magnitude adder
module sign_mag_add #(parameter N=4)
							(input  logic [N-1:0] a, b,
							 output logic [N-1:0] sum);
	
	// signal declaration
	logic [N-2:0]  mag_a, mag_b, mag_sum, max, min;
	logic sign_a, sign_b, sign_sum;
	
	// body
	always_comb
	begin
		// separate magnitude and sign
		mag_a = a[N-2:0];
		mag_b = b[N-2:0];
		sign_a = a[N-1];
		sign_b = b[N-1];
		// sort according to magnitude
		if (mag_a > mag_b)
			begin
				max = mag_a;
				min = mag_b;
				sign_sum = sign_a;
			end
		else
			begin
				max = mag_b;
				min = mag_a;
				sign_sum = sign_b;
			end
		// add/sub magnitude
		if (sign_a==sign_b)
			mag_sum = max + min;
		else
			mag_sum = max - min;
		// form output
		sum = {sign_sum, mag_sum};
	end  // always_comb
	
endmodule  // sign_mag_add


/* Testbench for Homework 2 Problem 4 */
module sign_mag_testbench ();

	// for you to implement BOTH sign_mag_add and sync_rom
	logic [3:0] a, b, sum;
	logic [7:0] addr;
	logic [3:0] data;
	logic clk;
	
	sign_mag_add #(4) dut (.*);
	sync_rom dut2 (.*);

	assign addr = {a, b};
	
	parameter CLOCK_PERIOD = 100;
	initial begin
		clk <= 0;
		forever #(CLOCK_PERIOD / 2) clk <= ~clk;
	end

	initial begin
	
//		// for you to implement
		@(posedge clk) a = 4'b0110; b = 4'b0000;  // pos + 0
		@(posedge clk);
		@(posedge clk) a = 4'b0110; b = 4'b1100;  // pos + neg valid
		@(posedge clk);
		@(posedge clk) a = 4'b0110; b = 4'b0001;  // pos + pos valid
		@(posedge clk);
		@(posedge clk) a = 4'b1110; b = 4'b1001;  // neg + neg valid
		@(posedge clk);

		@(posedge clk) a = 4'b1110; b = 4'b0110;  // pos + neg = 0
		@(posedge clk);
		@(posedge clk) a = 4'b1110; b = 4'b1111;  // pos + neg < 0
		@(posedge clk);
		@(posedge clk) a = 4'b0110; b = 4'b0110;  // pos + pos overflow
		@(posedge clk);
		@(posedge clk) a = 4'b1110; b = 4'b1110;  // neg + neg overflow
		@(posedge clk);
		@(posedge clk);
		
		$stop;
	end  // initial
	
endmodule  // sign_mag_testbench
