module DE1_SoC (
	);
	
	
	
endmodule  // DE1_SoC
